`timescale 1ns / 1ps

module tb_TensorUnit();
    parameter   D_WIDTH = 32,
                M_SIZE  = 4;
    reg aclk;
    reg aresetn;
    
    reg  [(D_WIDTH) * (M_SIZE) * (M_SIZE) - 1:0]  i_matrix;
    reg  [(D_WIDTH) * (M_SIZE)            - 1:0]  i_vector;
    wire [(D_WIDTH) * (M_SIZE)            - 1:0]  o_result;
    
    reg  [(D_WIDTH) * (M_SIZE) * (M_SIZE) - 1:0]  MATRIX_2X2;
    reg  [(D_WIDTH) * (M_SIZE) * (M_SIZE) - 1:0]  MATRIX_3X3;
    reg  [(D_WIDTH) * (M_SIZE) * (M_SIZE) - 1:0]  MATRIX_4X4;
    reg  [(D_WIDTH) * (M_SIZE) * (M_SIZE) - 1:0]  MATRIX_10X10;
    
    reg  [(D_WIDTH) * (M_SIZE)            - 1:0]  VECTOR_2X1;
    reg  [(D_WIDTH) * (M_SIZE)            - 1:0]  VECTOR_3X1;
    reg  [(D_WIDTH) * (M_SIZE)            - 1:0]  VECTOR_4X1;
    reg  [(D_WIDTH) * (M_SIZE)            - 1:0]  VECTOR_10X1;
    
    
    
    reg i_matrix_is_valid;
    reg i_vector_is_valid;
    reg i_receiver_ready_for_result;
    wire o_ready_to_accept_matrix;
    wire o_ready_to_accept_vector;
    wire o_result_is_valid;
    wire o_this_is_the_last_result;
    reg [31:0] temp;
    
    
    
    
    
    initial begin
        aclk = 0;
        forever aclk = #5 ~aclk;
    end
    
    TensorUnit #(.D_WIDTH(D_WIDTH), .M_SIZE(M_SIZE)) TensorUnit_Inst (
        .aclk                       ( aclk                          ),
        .aresetn                    ( aresetn                       ), 
        .i_matrix_is_valid          ( i_matrix_is_valid             ),
        .i_vector_is_valid          ( i_vector_is_valid             ),
        .i_receiver_ready_for_result( i_receiver_ready_for_result   ),
        .o_ready_to_accept_matrix   ( o_ready_to_accept_matrix      ),
        .o_ready_to_accept_vector   ( o_ready_to_accept_vector      ),
        .o_result_is_valid          ( o_result_is_valid             ),
        .i_matrix                   ( i_matrix                      ),
        .i_vector                   ( i_vector                      ),
        .o_result                   ( o_result                      ),
        .o_this_is_the_last_result  ( o_this_is_the_last_result     )
    );
    
    initial begin
        MATRIX_2X2 = { {32'b00111111_100000000_000000000_000000}, {32'b01000000_00000000_00000000_00000000}, // 2, 1
                        {32'b01000000_10000000_00000000_00000000}, {32'b01000001_00000000_00000000_00000000}}; // 4, 8 = 12
         VECTOR_2X1 = { {32'b01000000_01000000_00000000_00000000}, {32'b01000000_10100000_00000000_00000000}}; // 3, 5     
         
         MATRIX_3X3 = { {32'b01000000100110111010100110000010},{32'b01000000110001000001011100110001},{32'b00111111111010010110111111111011},
                        {32'b01000001000100101011010111101001},{32'b01000001000111110110011010111000},{32'b01000000110100110100011101001101},
                        {32'b01000000101110011000000010011101},{32'b01000001000101111111011001011110},{32'b01000000101111001011110010000011}};
         VECTOR_3X1 = { {32'b01000000110010011010010110101011},{32'b01000001000001110011011001100000},{32'b01000000000110111000101011110100}};
         
         
         MATRIX_4X4 = { {32'b01000000100110111010100110000010},{32'b01000000110001000001011100110001},{32'b00111111111010010110111111111011},{32'b01000000111111011101110100110000},
                        {32'b01000001000100101011010111101001},{32'b01000001000111110110011010111000},{32'b01000000110100110100011101001101},{32'b01000000100100000010111000100001},
                        {32'b01000000101110011000000010011101},{32'b01000001000101111111011001011110},{32'b01000000101111001011110010000011},{32'b01000001000011110011010011001011},
                        {32'b01000001000001111110101011110001},{32'b01000001000000011101110001001111},{32'b01000000001100000110011111100100},{32'b01000000111000011011000011010000}};
         VECTOR_4X1 = { {32'b01000000110010011010010110101011},{32'b01000001000001110011011001100000},{32'b01000000000110111000101011110100},{32'b01000000111010100001001110011000}};


         MATRIX_10X10 = { {32'b01000001000001110001101110000100},{32'b01000000111100101000101110011111}, {32'b01000000100001101001010100111001},{32'b01000000001001011011010011101011},{32'b01000000101000111001101110100000},{32'b01000000100000011001010000110100},{32'b01000000111110101101000011000111},{32'b01000000010000100001111011000001},{32'b01000000100110001000001011010010},{32'b01000000101110101010111010101000},
                          {32'b01000001000100010100110001001101},{32'b01000000101000010111111111110010}, {32'b01000000001101000110000001001111},{32'b01000000111100011101101101111010},{32'b01000000110001011110000011001001},{32'b01000000001000000101001011110101},{32'b01000001000100011000111100110100},{32'b01000001000111010011111011100100},{32'b01000001000000011010001001111111},{32'b01000001000100000101100010110111},
                          {32'b01000000010001100111111010010011},{32'b01000000111010011000101111010001}, {32'b01000001000011111101000001101010},{32'b01000000110110101101111111110110},{32'b01000000100101110001010111101110},{32'b00111111100000001110010111000101},{32'b01000000100010101110111101011011},{32'b01000000110000110111101111011100},{32'b01000001000100100001010011101110},{32'b01000001000110101010100000110010},
                          {32'b01000000100110001010010010100100},{32'b01000001000010100111001100011000}, {32'b01000000001001101011011100001111},{32'b01000001000000001100110111110000},{32'b01000000101011111001010101110010},{32'b00111111100100011111100100101111},{32'b01000000111001100100111000110101},{32'b01000000011111110011111100111111},{32'b01000001000000111111100110100110},{32'b01000000110101011100111100011100},
                          {32'b00111100001110110011110101010001},{32'b01000000100111011111000111100110}, {32'b01000001000010101101000100000010},{32'b01000000000111000001101001011011},{32'b01000000010100000010000101111011},{32'b01000001000010110100011010000000},{32'b00111111111101001001000011011101},{32'b01000000101101011001101001111010},{32'b01000000000110001011011011010101},{32'b01000001000110101100111001110010},
                          {32'b01000001000000001000001000111011},{32'b01000000100011110101100110101010}, {32'b00111111111001101111100001111100},{32'b01000000010011001101010110111111},{32'b01000000101000101000101001111111},{32'b01000001000101010100000011011111},{32'b00111111100010111001100000010011},{32'b01000000101100000110011111010000},{32'b01000000111000100001100110000010},{32'b01000000101011110010111001011100},
                          {32'b01000001000000100101000010010000},{32'b01000000101011001110010000001000}, {32'b01000001000110100011011011010011},{32'b01000000110000010000010011110111},{32'b01000000101111000000100110010111},{32'b01000000100011100110010110000000},{32'b01000000101111101100111111010001},{32'b01000000011101100101011000110100},{32'b01000000101110000011010101010100},{32'b01000000001110011100111110010101},
                          {32'b00111111111100100110101111000000},{32'b00111111111011110000001110001000}, {32'b01000000110001000001011001100000},{32'b01000000110100100010000110001001},{32'b01000000100110000111110101101011},{32'b00111111111100101111100110100101},{32'b01000000111100100110111011101001},{32'b01000001000011000100100010000011},{32'b01000001000100111011110110101111},{32'b01000001000001101100101100101011},
                          {32'b01000001000011111011010100101011},{32'b01000001000100111011000101110100}, {32'b01000000101011001111110111110010},{32'b01000000011110100110110111110001},{32'b01000000111000011011000011010000},{32'b01000000001100000110011111100100},{32'b01000001000000011101110001001111},{32'b01000001000001111110101011110001},{32'b01000001000011110011010011001011},{32'b01000000101111001011110010000011},
                          {32'b01000001000101111111011001011110},{32'b01000000101110011000000010011101}, {32'b01000000100100000010111000100001},{32'b01000000110100110100011101001101},{32'b01000001000111110110011010111000},{32'b01000001000100101011010111101001},{32'b01000000111111011101110100110000},{32'b00111111111010010110111111111011},{32'b01000000110001000001011100110001},{32'b01000000100110111010100110000010}};
        
         VECTOR_10X1 = { {32'b01000000110010011010010110101011},{32'b01000001000001110011011001100000}, {32'b01000000000110111000101011110100},{32'b01000000111010100001001110011000},{32'b00111111100101011110111010010000},{32'b01000000000011010001100001000001},{32'b01000000111111100100010000111100},{32'b01000000010101001101001010111001},{32'b01000001000000101000101111001100},{32'b00111111100000001100011100010010}};
    end
    
    initial begin
        // initial signal conditions
        i_receiver_ready_for_result = 1'b0;
        i_matrix_is_valid           = 1'b0;
        i_vector_is_valid           = 1'b0;
        i_matrix = {(D_WIDTH*M_SIZE*M_SIZE){1'b0}};
        i_vector = {(D_WIDTH*M_SIZE       ){1'b0}};
        
        aresetn = 1'b1; #20 aresetn = 1'b0;
        
        #20 aresetn = 1'b1; #20;
        
        
        /*
         *  | 8  4 |     | 5 |   | 52 |
         *  | 2  1 |  x  | 3 | = | 13 |
         */
         
         i_matrix = MATRIX_4X4;
         i_vector = VECTOR_4X1;    

        
        #10;
        // Check the ready signal and assert the valid signals
        if ( o_ready_to_accept_matrix &  o_ready_to_accept_vector) begin
            $display("[*] Matrix and Vector Valid");
            i_matrix_is_valid = 1'b1;
            i_vector_is_valid = 1'b1;
        end else begin
            $display("[*] Matrix and Vector Invalid");
            i_matrix_is_valid = 1'b0;
            i_vector_is_valid = 1'b0;
        end
        
        /* DELAY    */    
        #60;
        // Assert that the receiver is ready to receive the data
        i_receiver_ready_for_result = 1'b1;
        
        #10;
        i_matrix_is_valid = 1'b0;
        i_vector_is_valid = 1'b0;
        
        #10;
        if (o_this_is_the_last_result) begin
            $display("Last result obtained");
            $display("o_result = %d", o_result);
        end
 
    end
endmodule