`timescale 1ns / 1ps

// Verilog-2005 does not allow two dimensional arrays in the input/output ports
// Therefore, we can do it with custom macros.
`include "preprocessors.v"

module TensorUnit #(parameter D_WIDTH=32, M_SIZE=2) (
    // SYSTEM SIGNALS
    input   aclk,
    input   aresetn,
    
    // AXI CONTROLS 
    input   i_matrix_is_valid,
    input   i_vector_is_valid,
    input   i_receiver_ready_for_result, // input to the accumulator
    //input   i_accumulator_waiting_for_data, // output from accumulator
    output  o_ready_to_accept_matrix,
    output  o_ready_to_accept_vector,
    output  o_result_is_valid,
    output  o_this_is_the_last_result,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   
    // DATA
    input  [(D_WIDTH) * (M_SIZE) * (M_SIZE) - 1:0]  i_matrix,
    input  [(D_WIDTH) * (M_SIZE)            - 1:0]  i_vector,
    
    output [(D_WIDTH) * (M_SIZE)            - 1:0]  o_result
);
    
    // Internal data registers and wires
    reg  [D_WIDTH-1:0] r_partial_matrix    [0:M_SIZE-1][0:M_SIZE-1];
    wire [D_WIDTH-1:0] w_partial    [0:M_SIZE-1][0:M_SIZE-1];    
    wire [D_WIDTH-1:0] wi_matrix    [0:M_SIZE-1][0:M_SIZE-1];
    wire [D_WIDTH-1:0] wi_vector    [0:M_SIZE-1];
    wire [D_WIDTH-1:0] wo_vector    [0:M_SIZE-1];
    wire [D_WIDTH-1:0] w_o_result   [0:M_SIZE-1];
    
    // Loop controls
    integer count_x, count_y;
    
    // Unpack the arrays : see the template
    `UNPACK_MATRIX(D_WIDTH, M_SIZE, wi_matrix, i_matrix)
    `UNPACK_VECTOR(D_WIDTH, M_SIZE, wi_vector, i_vector)
    
    
    // Internal interfacing signals for MATRIX_VECTOR_MULTIPLIER
    wire w_s_axis_partial_tvalid_all;
    wire w_m_axis_i_matrix_ready [0:M_SIZE-1][0:M_SIZE-1];
    wire w_m_axis_i_vector_ready [0:M_SIZE-1][0:M_SIZE-1];
    wire w_s_axis_partial_tvalid [0:M_SIZE-1][0:M_SIZE-1];
    
    // Internal interfacing signals for ACCUMULATOR
    
    /* Here, the following block multiplies all the matrix elements with the vector and stores the result in partial matrix */
    /* 
     * If M_SIZE = 3, then, by the end of this operation, we will have the following result.
     * NOTE: we still need to add the elements in each row.
     * a[i][j] x b[j] = partial_matrix[a[i][j]*b[i]]
     * 
     * | a[0][0] a[0][1] a[0][2] |     | b[0] |    | a[0][0]*b[0]   a[0][1]*b[1]   a[0][2]*b[2] |
     * | a[1][0] a[1][1] a[1][2] |  x  | b[1] | =  | a[1][0]*b[0]   a[1][1]*b[1]   a[1][2]*b[2] |
     * | a[2][0] a[2][1] a[2][2] |     | b[2] |    | a[2][0]*b[0]   a[2][1]*b[1]   a[2][2]*b[2] |
     */
     
    genvar row, element;
    generate
        for (row = 0; row < M_SIZE; row = row + 1) begin
            for (element = 0; element < M_SIZE; element = element + 1) begin
                // Instantiate the floating point ip
                fp_multiply_ab MATRIX_VECTOR_MULTIPLIER (
                    .aclk                   ( aclk                                  ),      // input wire aclk
                    .aresetn                ( aresetn                               ),      // input wire aresetn
                    .s_axis_a_tvalid        ( i_matrix_is_valid                     ),      // input wire s_axis_a_tvalid
                    .s_axis_a_tready        ( w_m_axis_i_matrix_ready[row][element] ),      // output wire s_axis_a_tready
                    .s_axis_a_tdata         ( wi_matrix[row][element]               ),      // input wire [31 : 0] s_axis_a_tdata
                    .s_axis_b_tvalid        ( i_vector_is_valid                     ),      // input wire s_axis_b_tvalid
                    .s_axis_b_tready        ( w_m_axis_i_vector_ready[row][element] ),      // output wire s_axis_b_tready
                    .s_axis_b_tdata         ( wi_vector[element]                    ),      // input wire [31 : 0] s_axis_b_tdata
                    .m_axis_result_tvalid   ( w_s_axis_partial_tvalid[row][element] ),      // output wire m_axis_result_tvalid
                    .m_axis_result_tready   ( w_accumulator_waiting_for_data[row]   ),      // accumulator is ready for input  /// LOOK OUT FOR THIS!
                    .m_axis_result_tdata    ( w_partial[row][element]               )       // output wire [31 : 0] m_axis_result_tdata
                );
                
                
            end
        end
    endgenerate
    
    assign o_ready_to_accept_matrix    = w_m_axis_i_matrix_ready[0][0];
    assign o_ready_to_accept_vector    = w_m_axis_i_vector_ready[0][0];
    assign w_s_axis_partial_tvalid_all = w_s_axis_partial_tvalid[0][0];
    
    
    /* If all of the partials are calculated, then assign it to a temporary memory */
    /* This is in case we need to pipeline the whole design. */
    always @(w_s_axis_partial_tvalid_all) begin
        if (w_s_axis_partial_tvalid_all) begin 
            for (count_x = 0; count_x < M_SIZE; count_x = count_x + 1)
                for (count_y = 0; count_y < M_SIZE; count_y = count_y + 1) begin
                    r_partial_matrix[count_x][count_y] = w_partial[count_x][count_y];
                end
        end  else begin
           r_partial_matrix[count_x][count_y] = 0;
        end
    end
    
    
    /* The first part is done, we begin the second stage of the calculation */
    
    
    reg r_external_receiver_ready,
        r_input_data_is_valid,
        r_last_input_to_accumulator;
        
    reg  [D_WIDTH-1:0]  r_matrix_row_element                    [0:M_SIZE-1];
    wire [D_WIDTH-1:0]  w_accumulated_row_sum                   [0:M_SIZE-1];
    
    wire                w_accumulator_waiting_for_data          [0:M_SIZE-1],
                        w_accumulator_result_is_valid           [0:M_SIZE-1],
                        w_last_result_before_accumulator_reset  [0:M_SIZE-1];
    
    
    /* We will need a state machine for shifting the values in to the accumulator */
    localparam  IDLE = 2'b00,
                LOAD = 2'b01,
                NEXT = 2'b10,
                NOP  = 2'b11;
    reg [1:0]   state;                
    reg [4:0]   row_idx, col_idx;
    
    
    always @ (posedge aclk or negedge aresetn) begin
        if (!aresetn) begin
            r_external_receiver_ready   <= 1'b0;
            r_input_data_is_valid       <= 1'b0;
            col_idx                     <= 0;
            state                       <= IDLE;
            
        end else begin
            
            if (w_s_axis_partial_tvalid_all) begin
            
                /* assert data is valid as all partials have been calculated */
                r_input_data_is_valid       <= 1'b1;
                r_external_receiver_ready   <= i_receiver_ready_for_result;
                
            end else begin
                r_input_data_is_valid       <= (!r_last_input_to_accumulator) ? r_input_data_is_valid : 1'b0;;
                r_external_receiver_ready   <= 1'b0;
            end
            
            /* control path: we now shift the elements of the partial matrix one by one to the input to the accumulator */
            case (state)
            
                IDLE:   state <= (r_input_data_is_valid) ? LOAD : IDLE;
                
                LOAD:   
                begin
                    if (col_idx < M_SIZE) state <= LOAD;
                    else                          state <= IDLE;                     
                    
                    if (o_this_is_the_last_result) state <= IDLE;
                    
                    col_idx         <= col_idx + 1;
                end
                
                default:state <= IDLE;
            endcase
            
        end
    end
    
    always @* begin
        for (row_idx = 0; row_idx < M_SIZE; row_idx = row_idx + 1) begin
            /* data path: we now shift the elements of the partial matrix one by one to the input to the accumulator */
            case (state)
                IDLE: begin
                      r_matrix_row_element[row_idx]   = {M_SIZE, {1'b0}};   
                      r_last_input_to_accumulator     = 1'b0;
                end       
                LOAD: begin
                        r_matrix_row_element[row_idx]       = (col_idx < M_SIZE) ? r_partial_matrix[row_idx][col_idx] : 0;
                        
                        if (col_idx == (M_SIZE - 1))  
                            r_last_input_to_accumulator     = 1'b1;
                        else
                            r_last_input_to_accumulator     = 1'b0;
                end
                default: r_matrix_row_element[row_idx]   = {M_SIZE, {1'b0}};
            endcase
        end
    end
    
    integer sum_idx;
    reg [D_WIDTH-1:0] temp_sum [0:M_SIZE-1];
    always @(posedge aclk or negedge aresetn) begin
        if (!aresetn) begin
            for (sum_idx = 0; sum_idx < M_SIZE; sum_idx = sum_idx + 1)
                temp_sum[sum_idx] <= 0;
        end else begin
            if (o_this_is_the_last_result)
            for (sum_idx = 0; sum_idx < M_SIZE; sum_idx = sum_idx + 1)
                temp_sum[sum_idx] <= w_accumulated_row_sum[sum_idx];
        end
    end
    
    genvar adder_row_idx;
    generate
        for (adder_row_idx = 0; adder_row_idx < M_SIZE; adder_row_idx = adder_row_idx + 1) begin                
              fp_accumulator_ai ACCUMULATE_PARTIAL_ROW_0 (
                  .aclk                 ( aclk                                                  ),
                  .aresetn              ( aresetn                                               ),
                  .s_axis_a_tvalid      ( r_input_data_is_valid                                 ),  // input wire : incoming data valid?
                  .s_axis_a_tready      ( w_accumulator_waiting_for_data[adder_row_idx]         ),  // output wire s_axis_a_tready
                  .s_axis_a_tdata       ( r_matrix_row_element[adder_row_idx]                   ),  // input wire [31 : 0] : elements from partial matrix
                  .s_axis_a_tlast       ( r_last_input_to_accumulator                           ),  // input wire s_axis_a_tlast
                  .m_axis_result_tvalid ( w_accumulator_result_is_valid[adder_row_idx]          ),  // output wire : is the output data valid?
                  .m_axis_result_tready ( i_receiver_ready_for_result                           ),  // input wire : this is master, slave is ready for accepting data
                  .m_axis_result_tdata  ( w_accumulated_row_sum[adder_row_idx]                  ),  // output wire [31 : 0] : row-wise sum available here
                  .m_axis_result_tlast  ( w_last_result_before_accumulator_reset[adder_row_idx] )   // output wire, last calculated data
                );
                
        end
    endgenerate

    assign o_this_is_the_last_result = w_last_result_before_accumulator_reset[0];
    assign o_result_is_valid         = w_accumulator_result_is_valid[0];
    
    `PACK_VECTOR(D_WIDTH, M_SIZE, o_result, temp_sum)
endmodule

